LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY decod_4_16 IS
	PORT( a: in std_logic_vector(3 downto 0);
			s: out std_logic_vector(15 downto 0)
	);

END decod_4_16;

architecture arq_decod_4_16 of decod_4_16 is
	begin
		WITH a SELECT
			s <=
				"0000000000000001" WHEN "0000",
				"0000000000000010" WHEN "0001",
				"0000000000000100" WHEN "0010",
				"0000000000001000" WHEN "0011",
				"0000000000010000" WHEN "0100",
				"0000000000100000" WHEN "0101",
				"0000000001000000" WHEN "0110",
				"0000000010000000" WHEN "0111",
				"0000000100000000" WHEN "1000",
				"0000001000000000" WHEN "1001",
				"0000010000000000" WHEN "1010",
				"0000100000000000" WHEN "1011",
				"0001000000000000" WHEN "1100",
				"0010000000000000" WHEN "1101",
				"0100000000000000" WHEN "1110",
				"1000000000000000" WHEN "1111",
				"----------------" WHEN others;

end arq_decod_4_16;